LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;
use IEEE.STD_LOGIC_arith.all;
use IEEE.std_logic_textio.all;
use IEEE.numeric_bit.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_signed.all;
use IEEE.std_logic_unsigned.all;
use IEEE.math_real.all;
use IEEE.math_complex.all;

ENTITY tdes_tb IS
END tdes_tb;

ARCHITECTURE tdes_tb_behav OF tdes_tb IS

	-- Importação de componente
	COMPONENT tdes port (
		clock          : IN std_logic;
		reset          : In std_logic;
		text64         : IN std_logic_vector(0 TO 63);
		key192         : IN std_logic_vector(0 TO 191);
		done           : OUT std_logic;
		textOut64      : OUT std_logic_vector(0 TO 63)
		);
	END COMPONENT;

	signal sig_clock        : std_logic;
	signal sig_reset        : std_logic;
	signal sig_text64       : std_logic_vector(0 TO 63);
	signal sig_key          : std_logic_vector(0 TO 63);
	signal sig_done         : std_logic;
	signal sig_textOut64    : std_logic_vector(0 TO 63);
BEGIN
	-- Mapeamento de portas
	UUT_des_box: tdes PORT MAP(
		clock     => sig_clock    ,
		reset     => sig_reset    ,
		text64    => x"726f646f6c666f31"   ,
		key192    => x"133457799BBCDFF1133457799BBCDFF1133457799BBCDFF1",
		--text64    => x"13f666c6f646f627"   ,
		--key192    => x"1ffdcbb9977543311ffdcbb9977543311ffdcbb997754331",
		done      => sig_done     ,
		textOut64 => sig_textOut64
	);

	processClk: Process 
	BEGIN
		sig_clock <= '0';
		wait for 1 ns;
		sig_clock <= '1';
		wait for 1 ns;
	END PROCESS;

	-- Processo responsavel pela variação no dado de entrada
	signal_dadoA: PROCESS
	BEGIN
		--0123456789ABCDEF
		--key-133457799BBCDFF1

		sig_reset <= '1';
		wait for 2 ns;
		sig_reset <= '0';
		wait for 600000 ns;

	END PROCESS;

END ARCHITECTURE tdes_tb_behav;